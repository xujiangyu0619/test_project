module rst_gen # 
(
    parameter   CH  = 1
)
(
    input               clk,
    input       [7:0]   dat,
    input       [7:0]   key,
    output      [7:0]   led,

    output      [7:0]   line 
);


reg     [7:0]   reg_1;
wire    [7:0]   wire_1;


endmodule
