// pll.v module
module pll
();

endmodule
