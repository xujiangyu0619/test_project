module top 
(
    input       clk     ,
    input       rst_n   ,

    output      led     
);




endmodule
