// clock generate module
module clk_gen
(
    input clk,
    input rst_n,

    output led
);

    
endmodule
