// clock generate module
module clk_gen
(
    input clk,
    input rst_n,

    output led
);

reg     [7:0]   cnt;
    
endmodule
